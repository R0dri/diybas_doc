* AC Analysis, 600E-3 highPass, 4th order Butterworth, 2 stages using AD8602

*******************
* Supply Voltages *
*******************
VP VCCG 0 5
VR VGND 0 0
VM VEEG 0 -5


******************
* Import Signals *
******************
* Vtest testi 0 PWL (file=filters.txt)
Vin0 signal 0 PWL (file=signals/samplegit/data1/data0_1.csv)
*Vin IN     0 AC 1 PWL (file=signals/simulated/signals_src.txt)
Vcm1 VCM1   0 PWL (file=signals/simulated/signals_vcm.txt)
Vcm2 VCM2   0 PWL (file=signals/simulated/signals_vcm2.txt)
*XM VCM1 VCM2  VCCG VEEG VGND HPfilter

Vhp  HP     0 PWL (file=filters_hp.txt)
*Vina IA     0 PWL (file=filters_ina.txt)

Vin in 0 AC 1 DC 0 SIN(0 0 100)
***********
* Modulos *
***********
*R1 IN 1 1k
*R2 IN 2 1k
*R3 1 OUT_Ib 2k
*R4 2 VGND 2k
*    in  out            +5v   0v  2.5v
XH   IN      OUT_HP            VCCG VEEG VGND HPfilter
XC   OUT_HP  OUT_Ia        GND VCCG VEEG VGND INA
*XI   1      OUT_Ib       2 VCCG VEEG VGND INA
*XN   OUT_Ia  OUT_N             VCCG VEEG VGND Notch_50
XA   OUT_Ia   OUT              VCCG VEEG VGND LPfilter
* XR  VCM  REF    VCCG VEEG REF_BUFFER
* xd  ref   vdrl   vccg veeg vgnd drl



*** Conditions ***
*.TEMP 27
*.OPTIONS CHGTOL=10F ITL1=1000 ITL2=40 ITL4=20 TRTOL=14
*.OPTIONS numdgt=7 plotwinsize=0
*** Type ***
.AC DEC 100 16E-4 10E6
* .TRAN 50us
*.TRAN 0s 0.1s 0s 0.1ms
* .NOISE V(OUT) VNOISE DEC 100 16E-3 10E3
*.PWL IN

* .PROBE V(REF) V(VDRL)
* .PROBE V(v50) V(vdc) V(vnoise)
* .PROBE V(vcm) V(base) V(artf)

.PROBE V(out_hp) V(out_lp) V(out_ia) V(out_ib) V(out_n)
.PROBE V(vcm1) V(IN) v(signal) V(vcm2) V(hp)
.PROBE V(out)



******************
* Modules import *
******************
.lib modules.lib



